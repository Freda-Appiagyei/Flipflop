----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    14:28:52 07/08/2021 
-- Design Name: 
-- Module Name:    dflipflop - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity dflipflop is
port(
CLK ,D ,iload: IN STD_LOGIC;
Q      :OUT STD_LOGIC
);
end dflipflop;

architecture Behavioral of dflipflop is
begin
  process(CLK)
    begin
	 if (rising_edge(clk)) then 
	    if (iload='1')then
	     Q<=D;    
	    end if;
	 end if;
	 end process;
end Behavioral;

